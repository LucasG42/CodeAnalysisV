[translated]
module main

fn main() {
	C.printf(c'Hello World\n')
}
